@@ -0,0 +1,9 @@
<svg width="35" height="35" viewBox="0 0 35 35" fill="none" xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink">
<circle cx="17.5" cy="17.5" r="17.5" fill="url(#pattern0)"/>
<defs>
<pattern id="pattern0" patternContentUnits="objectBoundingBox" width="1" height="1">
<use xlink:href="#image0_685_262" transform="scale(0.00588235)"/>
</pattern>
<image id="image0_685_262" width="170" height="170" xlink:href="data:image/png;base64,iVBORw0KGgoAAAANSUhEUgAAAKoAAACqCAYAAAA9dtSCAAAAAXNSR0IArs4c6QAAHUhJREFUeF7tXQl4VNXZ/s6dLEwAV1yqggFcUBZBBDcURUWtqNUKPypV/1rRSk2FmLk3PPp3/LFmZkJE0aqg9Xcpri21rVpwS1GQtiKoIIqCiWtdaAUVhpDM/f7nHTMYkrkzc5eZe+7kfs+TxyVn+c533pxz7rcK8imjBOrr6/duaWmpLC8vr0wkEpVCiL5E1EcIgZ+9dF3fk4h6ZhqEmbcKIf4thNjIzF8y80Yi+piImoUQyZ9QKPSZvxXGEhC+cL6TQDgcLgkGg8OZeWQgEBim6/oQIhpKRLsXSEabiWgNEa3GTyKRWNXc3Lxi/vz5rQWaX+ppui1QH3/88UBTU9MoIcQ4Zj6BiI4not6S7dYWIcRyZn6JmRu3bdv293A43CYZjwVhp1sBNRaL7cvMZzLzGUKIU4loj4JI2blJNjPz80S0uKys7JkZM2Z84tzQco9U9ECNxWIDmfknzDxRCHG43NthjjtmXiuEeEIIsSAUCr1nrre3WhclUKdOnVo6cODAs4noCiI6jYgC3toW09zqRNTIzPdWVFT8saqqqsX0CJJ3KCqgzp49+8DW1tYrFUX5byLaV3LZ54s9aBQeEELMK6ZTthiAKiKRyARFUaqY+RQiKoY1OQXiZcwc1TTtKSJipwZ1YxxPb2osFpug6/r1Qoij3RCeh+ZcJYT4dSgUWuhVwHoRqKKuru4CRVF+RUSDPQQWGVh9WwgRqaysXDBp0qSEDAzlyoOngDp79uyRuq7Padd75rpGv10nCQghXg0EAtdWV1e/4hXheAKo+EhKJBJ3ENEErwjWI3w+VVZW9svp06e/Lzu/UgM1HA4rFRUV05h5FhHtKrswPcrfFl3Xb2xpaZkjs9VLWqDW1dWNUhTlXiIa5lEAeI3t90pKSq6srq5ulJFx6YDa7hxyPRHVElGZjEIrYp7aFEWZU15efoNsRgOpgBqNRg8looeJ6MgiBoMXlgbtwEWhUOh1WZiVBqj19fUXJRKJu4QQu8ginBQfPXr0oB/84AdUUlJCGzdupK+++soWi71796Z99tmHmJk+//xz+vbbb22Nl6fO8Ny6NhQK4fnlOrkO1Hnz5lVs2rRpPhFd7Lo00jBw6KGH0oABA0hRlORvAa6PPvqIVq+G26h5wlgYs+N4H3zwAa1duzY5tmzEzH8ioks1TYO/rGvkKlBnzZrVv6ysDNaS4a5JIMPEw4YNo7594dDflV577TX67DNzTvm77LILHX/88TtA2nHUTz/9lFatWiWjGMDTukAgcP5111231i0GXQPqzTfffGwgEABIpXQeqayspMGDjQ1fuLJXrFhhat+GDh1K/fr1M+zz3nvv0bvvvmtqzAI2/g8RTVJV9YUCzrljKleAGo1Gf0JEePtI+VVfVlZGJ510EpWWlhruCd6q//jHP0zt2fDhw2n//fc37JNIJGjp0qWyvlnBN8yu16qqCuNLQanQQBXRaBQ2+v+R2cvp8MMPp/79+2fcCCunH05TnKqZSPInQIr1ufF4fHo4HIYfbEGokECFO94cIcQvC7Iyi5MIIejUU08lnKpGhK/0ZcuWUVub+fClE044gfBWNSKcqs8//7ylsS0u2Wq3/+vfv/8VhXJuKQhQ2z3uHySiyValUqh+ABHAZERff/118srfvn27JZYCgQAdffTRtPvuxsGtePviDewBerq0tHTijBkz4vnmNe9AbQfpQ0T0X/lejBPjQ3102GGHpR0K6iOcpJs329PUQC978sknp/36x8Tvv/8+vf32204spxBjFASseQUqQDpgwAAEn51bCIk5MQdACrCmo5aWluS17ASdeOKJBMV/Ovrkk0/o9delMQplXa4Q4sWSkpIJ+TxZ8wZU2Ox79OjxqBDix1lXKlEDqKSgmkpHW7Zsob/97W+OcAt96m677ZZ2LI98UO3EOzM/W1FRcU6+fATyBVQRi8XuYuYrHdnVAg6S6UTFu/S5555zhBtc/RUVFUVxoqYWIYR4ZOvWrVPyoQ3IC1BjsdgsZoYHlOfogAMOoCOOOMKQ78bGRtq6dautdcFn4LTTTjN8o0LpD/WXF4mZb9c0rcpp3h0HajQavZSI7nea0UKN16tXLxo7dqzhdM3NzfTWW2/ZYmfgwIE0aNAgwzGgVYBBwaskhKgKhUK3O8m/o0BtaGg4rq2tDSa2Hk4yWcixoEfFaWdkldq2bRu9+OKLthxIxowZQ7vumj5gQdd1evbZZwn6VA8TErudpaqqM+8kJ61D7Q4mMH57LZ9TFzzg6scTwIisOKSkxsqmp4UL4SuveCbmLtPf0jeBQOAYpxxZHDlRb7nllmBrayukK6UXlNmTCcr44447zrDbF198Qa+++qrZYZPts/0RrFmzhuD2VyS0LhgMjq6qqvra7nocAWpdXd2DiqLA0aRoCE4pPXumz8/b2tqavJ6t0Lhx4ygYDKbtinGhVZDRL9XKWtEH/qyapp1nN/GFbaBGo1E4PP/O6kJk7Qfn5oMOOsiQPVioNm3aZIp9WKQAVLyD0xEcst98801TY3qhMTNfrWnaXXZ4tQXUhoaGQ9ra2lZmSw1uh0G3+uI0xalqRPjyhwbADO277740cuRIwy7Lly+n//wHbp9FRy3MfLSmaW9YXZlloLbb8PEuPcrq5LL3Gz9+vOHX/4YNG+idd94xtQS4DsKFMB3ha3/RokVFde13XCdyuZaVlR1l1cxqGaixWGwmM//a1E55rHEm69GHH35oOm4q03PCSauXrGJWFKW+pqYmZIU/S0Ctq6sboSjKP4moxMqkXumT6cOnqakpGZBnhvDmBVjTkZ0PNDM8uNxWZ+axmqYtNcuHaaC2X/kAaVGooowEBoU/HKhT0aKd261bt47Wr19vSt7ZPPzh8ALHlyKndfF4fHg4HN5mZp2mgRqNRq8lojlmJvFi20zvSawHelToU81QNmU/gI8/gGInIcSvQqHQ/5pZpymg3nTTTX1LS0shyfSKQDMzS9wWYSjwFy0vLzf88LFq5jz99NOTiSyMrn+cqlajByQWaWfWtpeUlAytrq7OOeTWFFCj0SicTeB0UtR0zDHH0J57oiBfeoIKCaokKzRq1Cjae++9DbsiegCRqN2AnlRVFYaAnChnoLZn1/s7EX2XMqRIab/99qMRI0ZkXB287+GFb4X22msvGj16dMau+EjDx1o3oPG5Oq7kDNRoNIoYDBRzKGoCSAFWI8LHzpIlS2zpOzN5T2HeL7/8kv75T3yvFj2tUFUVf7VZcxnlBNRYLDaemRcXvdiIKNu1v3LlSvrXv/5lSxR4VmAeI0Kk68svv2xrDq901nV9Um1t7RPZ+M0FqEgagT/vorVAdRQSrmVcz0bkRDxTprgszFtErn7Z8Iebae2AAQOGZcsPkBWoKJHDzH/JOmORNIDnPTzwjQimTlz9VsNRoFGAIQHx/UZkxerlcfFPUVV1QaY1ZAVqJBJZJoQwds70uIQ6sw8PJ4SiGKmQ0N6Ol1O2dEEeyD+Vjx1fo6oqUuAbvlUzAjUSiYwRQnSPx1IH8cPL6cgjjzR0x0M4ygsvWEtql8nPFX6o8MoqIsfpnEHNzBM0TXvaqEM2oC4UQuSs68qZKw80BFCRZdqIcP2bzRSdzR/VSoZAD4gyJxaZuVHTtHGmgVpXV1epKAqM2cVemTmtbLKZO+HgjCeAGcrmj2rFLGtmfsnbsqIow2tqatJ6jhueqNFodDYRVUu+uLyy57Q/aibvKbxNFy9ebEs/m1dhFGBwZr5P07TL002VFqjhcLhHMBj8mIiM7YgFYNztKTL5o+IdiUA8M5RJo+BkXiszPEnWNl5WVrbf9OnTu8T4pAUqKpToup5RXSDZAvPCzimnnEJ4V6YjK/6ohxxyCB188MFpx+sOjtM5btI0VVXv7Nw2LVBjsdgLzGz4sM1xQk83g54Tnk5GgXhIC4n0kGbowAMPpCFDhqTtgi9+JLaARqE7kxDitVAo1MW41AWot956a7+WlhZErWXVsRazQLM5p1hJtpvNdGolYLAY9yAQCAzunLiiCxi7i2N0tg1GVug+ffqkbWY17Q5OZ5zSRlap7mQ6zSL/G1VVDXds0wWo3c0SlU5gMHPifWoUhmLHZzRTXlT8ASBboH/9i3dCodBOab93Amo4HN4vGAxCOVjUPqfZTtNsySesvE9Tc2Z6p6KNx9KiZxOl5d8nEonDZs6cuSMefSegRqPRq4jIVkYLy5xJ1BG2fqSfTEd2q5bg2kfQoJEvgZNZrSUSqRVWNFVVo6mOnYGKupfnWBm1WPogTgrXvtHXvpWKfZ1lk805u5tEo2aDzBJVVXekqtkB1Llz55bH4/F/F2N6nmwS6fj7Qpg599hjDzr22GMN2bIT6mJmrZK3bSsrK9srpfzfAdSGhoaT29raXpSc+byzl0kp76SZM5N51ooxIe+CcWeC81RVfRJT7wBqNBpFnPUN7vAjz6yZCuvCWwpeU05QMZXvcUIeBmPMVVU1WemxI1C7RfBeNqHCcoQv83TkJFAzlZq045idbX1e+n1HK1USqKgJFQwG4QiQPnOtl1Znk9dM5Xtw9SPRrt38+tnqBFhxeLG5bFm7t8Xj8d3D4fC3SaDGYrHhzLxKVm4LyRecpeE0bURWqkp3HitbVRQrvq6FlFEh5yopKRlXXV3dmALqz5j5nkIyIOtcSI6GqihG6ilYj6DwN5vEN7VelK+EQcHI6gXnFFin4vG818GVdQt24kvX9VBtbW19EqjRaPQ2InK8iJUnJJGGSRSayFT9GWBCSh/Y5s0QSvbAhGr0R4Cx7JhnzfDilba6rj9UW1t7SepEbWRm4zzgXlmVQ3xm06ViGivx/dkqomBcX4e68yYqivJGTU3N8NSJCkW/5+tDOYTT5DCZvKfweytpd4466ijaZ599DNm0k3zNybVLNlbLhg0beovZs2f3SSQSX0rGnOvswLMfTwCjUjtWcvhncnZBKAqy+HV3z6l0G6/r+sGiPUtft8jIZRb9cExBip/OYEWWFIAK6czNEBxSoOjvXFUa4ET9U7Ph12bm9nJbIcTpor6+fpKu6495eSH55B2+qdCtpvKl4nqGJ75ZkKZ4hFYB2VKcGi+fa5dlbCHElSISiYSEEDvcqWRhzufDl0BKArqu1wGoc4UQ1/hi8SUgqwSEEL9DSslHiGiyrEz6fPkSIKLFACqqz57mi8OXgMQSWAGgopZp5qT1Eq/AZ61bSKAZQEUMf3q/tm4hA3+RskuAmb8GUD8nIuN6MrKvwuevO0igDUCFZ8Vu3WG1/hq9KwEAdWuxV+Lz7vb4nKckAKC2dddkvT4MvCMBADVRiMwoSLgAj6TKykpCNmc4fcD2Dd/MTP6ZVkQJ52af7EkAfgd33323vUEc7J33qx8x7EgMhhCPTJVGHFyTP5QDEkDGlt/85jcOjOTMEAAqgvp2dWa470dBxpFzzjknGdFpFHbh9Jz+eM5JQEagOq6ewvUOkBpla3ZOnP5I+ZKAZEBNqqc+IKJ+Ti0YEZyoTOefok5J1J1xJAPqN46aUJEO5+yzz85YPtEdsfuzmpWAZEBNmlAdcUpBodspU6YQHIN98r4EJANq0inFETe/n//859S7d2/v75C/gqQEJANq0s3vdiL6hZ39gfoJocA+FY8EJAPqAtuhKNCNXnPNNf6VXzwYle5ETYai2A3uQ3bmkSNHFtk2+cuR6URNBvfZDZe+6qqrkiZRK4RITlSsQ4ocEMKSjUrbWBnf72NdApIBNRkuvbeu61D6mybEp0+bNs20rR5ZRpC+8eOPUW71e5o6dSrttpvvcWh6I/LQAbb+O+/sUukxDzPlNOSgVEqfjVYK9CKTyJgxY3KaKdUIuT8feyx9GoHLLruM9t7b9+E2JdA8NUYCuHvukSLBY0s8Hu9lK0naeeedZ1iENp38kGHkjjvuMBTtxRdfTPvvv3+eRO8Pa0YCX3zxBd1///1muuSlbeckaZbSTl5yySWEzHe5EhLULlq0yLD5BRdcQMgf6pP7EsCz7OGHH3adkc5pJy0l8v3pT39qWC803QqfeeaZjDXuJ0yYkEx345P7EkAFwd///veuM9I5kS/KTr9qlqvLL798Rw6lXPriA2rVKuMM7Hjv4t3rk/sSQJ7WZ5+Fdd11Gq+q6nPJN+rjjz8eaGpqQpCfKRvopZdemjHfZ+clrl+/nhYuXGi4cpQeh7+AT+5L4M9//jO9886OUqRuMdSmKMpuNTU1W2yV7zH7poTedN68eYSPKiOqrq72daluwaJ9Xui1b7vttqSO203qUr4HzFgpiIZaSZlKJaZb5KZNm+iBBx4gJK5NR9DL9uzZ7asIuYmPZDLhuXPnuspD++RdC6LFYrHxzLzYDHewSMEyZZYAUlwrK1eupLY2BMF+Tz/60Y8ILoM+uScB5IC999573WOgfWZd1yfV1tY+gf/ccfWHw+GyYDAIxb+pd+rVV19tWDLc9ZX6DFiSwJo1awgaGpepNRgM9qmqqvp6J6C2X/+my6CfccYZNGzYMJfX5E/vpAQefPBB+uyzz5wc0spY6cugtwMV9/hdZkZF6nC8K33PfjNSk7ctCrHdfjtclF0nTVXVHZnQd1z9YOvWW2/t19LSgux+O/3/bCwj4nTQoEHZmvm/94AEUDD4kUcQ9OEuMfMwTdNWp7joAshoNLqUiI43wyYiTvFW7Vztw8wYfls5JPD0008ni2m4TGtUVR3akYcuQI3FYtcws2ndRN++fWnSpEm+DtTlHbYzvSzXPjPfoGnaTdmAui8zw1E0YHbRsNP/8Ic/9GP6zQpOkvarV6+mv/71r65zI4Q4KBQKbcgIVPwyFou9wMzjrHA8atQoGjt2rA9WK8JzsQ8SyyEpmgRF2VaqqtoltintR5PdOCqcrOPHjydoBHzyhgSgjoJaym1i5qmapnXx2E4L1Hbl/0d2UqYjxv/cc89NZvFzOq2k28Istvlxmj700EP0+eeWIpKcFMc38Xh8v3A4/G3nQQ3VULFYrJ6Zr7PLBT6ykIsKZlE/H5Vdaean/yeffEILFizIz+DmRv2tqqo/S9fFEKgNDQ2HtLW1ve1Ukl+csPA1xQmLf0daSh+45nYxH61xmt53330E+77bpOv66Nra2rR+0RkV+5FIZKEQ4jy3F+AbFPK3A01NTfTEE0m/D1eJmRs1TTP8gM8G1DFCiJddXQHMZEIkzbS+QcHZnYBfMEKiZUglz8wTNE172miFWU2lsVhsBTO7ngoFji9wgPHJGQnAORo6U3hKSUDvxePxQeFw2LD4Qi5AncDMf5FgMTRx4kTq37+/DKx4nofm5maEIMmyjimqqmb8mssKVKwkGo0uJ6Jj3F4V0v3AUduPALC3EzCVIiTI7VCT9lWsjsfjwzOdpmiXE1CteP/bE6VxbwQATp482a+wYlHAiKh49NFH6dNPP7U4grPdOnrxZxo5J6BigEgkskwIIUUs89ChQ5PvVd+QYA40eJc+//zzGUPWzY1ou/WaeDx+RLbTNOcTFQ1jsdhwZl5hxVnF9nLSDHDWWWfR4MGD8zF00Y65bt06+tOfEMQhBbEQ4oRQKLQsF25yPlHb36rzieiKXAYuRBsEAqLAhU/ZJSDZxxNuwydCodCk7Jx/18IUUNtTVK6TqRr1hRdeSDDT+mQsAVnySHXgcEtra+th119/PfxJciJTQMWI9fX1M3Rdb8hp9AI0wjsV2VVgmvWpqwSQlQ95FFLJkiWR0Y2qqobN8GIaqOFwWAkGgy+ZDVcxw5SVttAE9OvnWF03KyxI1wdf9sjIJ4PlqYNwVsXj8dHhcHjnhA5ZpGcaqBjv5ptvHhQIBF4nonKZdgduhXizdndtAE5PxD1JEJvfGR4JXdePNXI8yYQlS0DFgJFI5NdCiJkyARW8wNSKAhjdNXwbelJk4ZPENLoTPBRFubOmpmaaFcxYBmo4HC5pfwIca2XifPbBxxVO1+7mxIICEcjCh5BnCenNYDA4uqqqKn3SsXxc/akx58yZM6ClpWWVEMJaWZQ8ShPXP9RXBx10UNE/BXDVI6Xnk08+KdtHU2qH48w8StM0y3HYlk/UFAeRSORKIcTdecScraFRURDBhsVakh2pPJcsWZJMOCcrpbJG2+HPNlAxeTQaReq3y+0wks++qC6IpwA8r4olqgBf8qgw89RTTxGcTGQlZn5c07TJRPRdMTGL5AhQw+Fwj4qKipdwvFvkoyDd9thjDzrzzDMJji1e1QzgmkcQHgAqQ/hIlo17Kx6PH5MuWM/shjsCVEx600039S0tLX2NiKRPbjpw4EA66aSTCMD1CmABUABz+fLltHbtWrP77Eb7zSUlJaOrq6vfdWJyx4AKZurq6k5VFAWJNUudYC7fY0A7cPLJJyeLsMn6JEgkEskUkI2NjdK45uWwL7qu6xfU1tb+MYe2OTVxFKiYMRKJTBZCoECR42PntCILjRAVe+KJJybfsDKotHB6fvPNN4TAu2XLlsmQvcSUVIUQVaFQyNHclXkBUywWm8XM15tanSSNAdYRI0YkfQcKGUkAcEIPihh7gHPjRiT/9h4x8+2aplU5zXlegAp/gIqKit8x84VOM1zI8XbffXcaMmQIHXDAAYR/d7L6NYCJKFC8O3FyvvHGG1J/veco96c2bNhw/vz581tzbJ9zs7wAFbOjdlVzc/ODzHxRztx4oCFKauJjDJlfevXqldTP4gdvXPykPs7wtoQKCf/EDyqNbN68OXlSfvjhh8nK2pJ5NNmVft5ACsbyBtQOYH2EmSfalYLfX2oJLIrH4+eGw+G8FabKK1Ah2ltuuSXY2tr6ByI6U2pR+8xZlcBLwWDw7FT1EquDZOuXd6B2OFnvZebLsjHk/947ElAUZeGWLVsuzOdJmpJGQYCaAmtTU9NviehS72yFz6mRBAoJ0ry/UdMtMhaL/ZKZ5+T7fexDLK8SQCjJjXbt92Y4LNiJ2pGpurq6iYqiIL1xDzPM+m1dl0CrEOLqUChU8PqTrgAV4m7PvvKYTBGtrsNAbga+1XX9EifNomaW6xpQwWQ0Gj1ACPEHZh5thmm/bcElsFrX9fNra2vXF3zm9gldBSp4mDt3bnk8Hr+DiNKmxHZLMP68OyTwWDwe/5kTrnp2ZOo6UFPMx2Kxacw823+32tlOR/tu13X9+traWuyJLadnJ7iSBqhYzKxZs/qXlZUhT6Z0AYNOCNtDY7wZCAQuvO6666RxfJUKqNjIdktWhIh+4VShCw8BxG1WcXL+Nh6PT3f7qu8sCOmAmmIwEokcoSjKPbKHt7iNLAfnfyuRSFwxc+ZMJG2WjqQFKiSFwmwVFRUaM9f6b9e8YQdv0Yby8vJZM2bMkDZKUGqgprYmHA7vV15eHlEUZYpv0XIOsLquP6QoykxVVVGkWWryBFBTEqyrqxunKArMr8Oklqr8zK1LJBIzZs6cifg2T5CngNoBsKcGAoGIDGWFPLHL7UwqivJGIpG4QdO0p2RQOZmRnSeBigUigqCpqekiJGpj5kFmFt0N224QQkTWr1//QD7CRAohT88CtaNwIpHIGEVRqpj5fFlqDBRi87LMAVXT08wc1TRtqQT82GKhKICakkAkEhkK7x7EacmYuM3WTuXeeQszPyaEuEtVVRQHKQoqKqCmdqS+vr6nruuTmfkKIcTRRbFT2RexkpnvraioWJDvsJDsrDjfoiiB2lFM7R5aP24PMESdrGJZM672V1BdZPv27QvNFG5wHkb5H7FYNi0nSTU0NByi6/oEXddR/fcEDxoRtgshluq6vhjvTzv5RnMSmESNuhVQO8p93rx5FV999dVYRVHG6bp+ghACFbRLJNobsJIQQqBWwku6rjdu27atUTYbfKHk1W2B2lnA4XC4VzAYPBa6WUVRhjHzECKC2qtQCd/amPldIcRqIlqdSCRW9erVa2kxvjetgNsHagapTZ06tXTgwIEDmLmSiCoVRalkZlRf6yOE6MPMSLG5JxH1zCL8rUT0byLayMxfKoqCxFIf67reTETN5eXlzZs3b95QiLBjKyCRoc//A9O+OVCSehUEAAAAAElFTkSuQmCC"/>
</defs>
</svg>
